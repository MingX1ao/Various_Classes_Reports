`timescale  1ns/1ns
module  tft_disp
(
    input   wire            tft_clk,    //���빤��ʱ��,Ƶ��33.3MHz
    input   wire            sys_rst_n,  //���븴λ�ź�,�͵�ƽ��Ч
    input   wire    [10:0]  pix_x,      //����TFT��Ч��ʾ�������ص�X������
    input   wire    [10:0]  pix_y,      //����TFT��Ч��ʾ�������ص�Y������

    output  reg     [23:0]  pix_data    //������ص�ɫ����Ϣ

);

//********************************************************************//
//****************** Parameter and Internal Signal *******************//
//********************************************************************//

parameter   H_VALID =   11'd800,   //����Ч����
            V_VALID =   11'd480;   //����Ч����

parameter   CHAR_B_H=   10'd272,   //�ַ���ʼX������
            CHAR_B_V=   10'd176;   //�ַ���ʼY������

parameter   CHAR_W  =   10'd256,   //�ַ����
            CHAR_H  =   10'd128;   //�ַ��߶�

parameter   BLACK   =   24'h000000,   //��ɫ
            GOLDEN  =   24'hFFD700;   //��ɫ

//wire  define
wire    [10:0]   char_x;   //�ַ���ʾX������
wire    [10:0]   char_y;   //�ַ���ʾY������

//reg   define
reg     [255:0] char    [127:0];   //�ַ�����

//********************************************************************//
//***************************** Main Code ****************************//
//********************************************************************//

//�ַ���ʾ����
assign  char_x  =   (((pix_x >= CHAR_B_H) && (pix_x < (CHAR_B_H + CHAR_W)))
                    && ((pix_y >= CHAR_B_V) && (pix_y < (CHAR_B_V + CHAR_H))))
                    ? (pix_x - CHAR_B_H) : 11'h3FF;
assign  char_y  =   (((pix_x >= CHAR_B_H) && (pix_x < (CHAR_B_H + CHAR_W)))
                    && ((pix_y >= CHAR_B_V) && (pix_y < (CHAR_B_V + CHAR_H))))
                    ? (pix_y - CHAR_B_V) : 11'h3FF;

//char:�ַ�����
always@(posedge tft_clk)
    begin
        char[0]     <=  256'h0000000000000000000000000000000000000000000000000000000000000000;
        char[1]     <=  256'h0000000000000000000000000000000000000000000000000000000000000000;
        char[2]     <=  256'h0000000000000000000000000000000000000000000000000000000000000000;
        char[3]     <=  256'h0000000000000000000000000000000000000000000000000000000000000000;
        char[4]     <=  256'h0000000000000000000000000000000000000000000000000000000000000000;
        char[5]     <=  256'h0000000000000000000000010000000000000000000000000000000000000000;
        char[6]     <=  256'h000000000000000000000001C000000000000000000000000000000000000000;
        char[7]     <=  256'h000000000000000000000001F000000000000000000000000000000000000000;
        char[8]     <=  256'h000000000070000000000001F800000000000000000000000000000000000000;
        char[9]     <=  256'h00000000007C000000000000FC00000000000000001E0000000000000007F000;
        char[10]     <=  256'h00003C00007E000000000000FC0000000000000001FF80000003C000007FF800;
        char[11]     <=  256'h00001F00007E000000000000F8000000000000003FFFE0000003F0180FFFF000;
        char[12]     <=  256'h00001F80007E000000000000780000000000001FFE07F0000001F81FFFFF0000;
        char[13]     <=  256'h00001F80007C000000000000780040000001FFFF8007F0000000FC0FFE000000;
        char[14]     <=  256'h00001F00007C0000000000007800F0000001FF83C007E00000007C0F00E00000;
        char[15]     <=  256'h00003F0000F80000000000007000F8000000F001E007C00000003C0F00F80000;
        char[16]     <=  256'h00003E0000F80000000000007000FC000000F001E007800000001C0F00F80000;
        char[17]     <=  256'h00003C0000F00000000000007001FE0000007001E00780000000000F00F80000;
        char[18]     <=  256'h00007C0001F00000000000007001FC0000007801E00780000000000F00F00000;
        char[19]     <=  256'h0000780001E00000000000007003F00000003801E00700000000000E00E00000;
        char[20]     <=  256'h0000F80001C00000000000007007E00000003801DF8F00000000000E00C00000;
        char[21]     <=  256'h0000F07C03C0380000000000700F800000001803FF0F00000078000E0181F000;
        char[22]     <=  256'h0000F0FE0380FE0000000000700F000000001C7FF80E0000007E000E018FF800;
        char[23]     <=  256'h0001E7FF0703FF80000000F0701E000000001C1DC00E0000003F001EC3FFFE00;
        char[24]     <=  256'h0001FFBF073F1FC0000007F87038000000000C01C00E0000003F001CFFF07E00;
        char[25]     <=  256'h0003C03E0FFC3FC000007FFC7070000000000C01C01C0000001F001CF0007E00;
        char[26]     <=  256'h000780381FF03F00001FFFF878E0000000000C01C01C0000000F001C70007C00;
        char[27]     <=  256'h0007803018007C00000FF0F07D80000000000E01C01C00000007001C70007C00;
        char[28]     <=  256'h000F006038007000000780F07F00000000000601C03800000000001C70007800;
        char[29]     <=  256'h000E00407000E000000001E07700000000000601DFF800000000003830FC7800;
        char[30]     <=  256'h001E380060008000000001E0738000000000060FFFF00000000004383FFE7800;
        char[31]     <=  256'h003C3E00CE000000000001E071C00000000007FFF0700000000008383FF07000;
        char[32]     <=  256'h00381E018F800000000003C070E00000000003F8006000000000183838007000;
        char[33]     <=  256'h00701E0007C00000000003C0707000000000030000000000000030703800F000;
        char[34]     <=  256'h00E01E0007C0000000000780707800000000000000003F00000030701800E000;
        char[35]     <=  256'h01C01C000780000000000780703C00000000000000001FE0000060701800E000;
        char[36]     <=  256'h03801C000780000000000F00701E00000000000000000FF00000E07018FFC000;
        char[37]     <=  256'h07001C000780000000000F00700F800000000001C00003F80000C0E01FFFC000;
        char[38]     <=  256'h06001C000780000000001E007007C00000060001F80001FC0001C0E018E08000;
        char[39]     <=  256'h00001C000780000000001C007007F00000060000FC0000FC000381E000700000;
        char[40]     <=  256'h000018000FC0000000003C007003FC0000060C007E00007C000381C000700000;
        char[41]     <=  256'h000018000FE00000000078007001FF80000F04003E00001C000781C000700000;
        char[42]     <=  256'h0000380C0F7000000000F0007000FFF0000F06001E010000000F03C000700000;
        char[43]     <=  256'h000038381E3800000001E00070007FFF001E06000E010000003F038080700000;
        char[44]     <=  256'h000038701E3800000001C000F0003FFFC01E030000018000007E07818070C000;
        char[45]     <=  256'h000039E01C1C000000038000F0001FFE003E03000000C000007E0701C070FC00;
        char[46]     <=  256'h00003BC03C0E000000070000F0000000003E03800000E000007C0F03C0707F00;
        char[47]     <=  256'h00007F80780F8000000E0000F0000000003C01C000007000007C0E0380703F80;
        char[48]     <=  256'h00007F007807C00000380000F0000000003C00E000007800007C1E0780701FC0;
        char[49]     <=  256'h0000FE00F003E00000700000F0000000003800F000007E0000781C0F80700FC0;
        char[50]     <=  256'h0001FC01E003F80000000040F00000000038007800007F000038380F007007C0;
        char[51]     <=  256'h0001F803C001FC000000003FF00000000030003E00007F800038700F007003E0;
        char[52]     <=  256'h0001F0078000FF800000001FF00000000000001FC007FF800010F00E007001C0;
        char[53]     <=  256'h0001E00F00007FF00000000FF00000000000000FFFFFFF000000E00C1FF00000;
        char[54]     <=  256'h0001C03C00007FFF00000007F000000000000003FFFFFC000001C0000FF00000;
        char[55]     <=  256'h000080F000003FFF80000003E0000000000000007FFFE0000003800007F00000;
        char[56]     <=  256'h0000008000001FFC00000003E00000000000000007FE00000006000003F00000;
        char[57]     <=  256'h000000000000000000000001C00000000000000000000000000C000001E00000;
        char[58]     <=  256'h000000000000000000000000C000000000000000000000000000000001E00000;
        char[59]     <=  256'h0000000000000000000000000000000000000000000000000000000000C00000;
        char[60]     <=  256'h0000000000000000000000000000000000000000000000000000000000000000;
        char[61]     <=  256'h0000000000000000000000000000000000000000000000000000000000000000;
        char[62]     <=  256'h0000000000000000000000000000000000000000000000000000000000000000;
        char[63]     <=  256'h0000000000000000000000000000000000000000000000000000000000000000;
        char[64]     <=  256'h0000000000000000000000000000000000000000000000000000000000000000;
        char[65]     <=  256'h0000000000000000000000000000000000000000000000000000000000000000;
        char[66]     <=  256'h0000000000000000000000000000000000000000000000000000000000000000;
        char[67]     <=  256'h0000000000000000000000000000000000000000000000000000000000000000;
        char[68]     <=  256'h0000000000000000000000000000000000000000000000000000000000000000;
        char[69]     <=  256'h0000000010000000000000000000000000000000180000000000000000000000;
        char[70]     <=  256'h000000003E0000000000000000000000000000003E0000000007000000000000;
        char[71]     <=  256'h000000007F8000000000000000000000000000001F0000000007C00000000000;
        char[72]     <=  256'h00000001FF8000000000000000000000000038001F0000000003E0003F000000;
        char[73]     <=  256'h00000007FC000000000000000078000000003E001F0000000003F0003FC00000;
        char[74]     <=  256'h0000003FC0000000000000003FFE000000001F001E0000000003F0001FE00000;
        char[75]     <=  256'h000000FE00C000000000007FFFFF800000000F001E0000000003F0000FE00000;
        char[76]     <=  256'h00000FE000F8000001E03FFF800FC00000000F001E7E00000001E00003E00000;
        char[77]     <=  256'h0000080000F8000000FFFFC0000FE000000007001FFF00000001E00001E00000;
        char[78]     <=  256'h0000001801F00000007FE0000007E0000000070FFFFF80000001E00000000000;
        char[79]     <=  256'h0000001C01E00000007800000007C00000001FFFFFFE00000001E00000000000;
        char[80]     <=  256'h0000301E03C00000007800000007C000003FFFF8380000000001E00000000000;
        char[81]     <=  256'h00003C0F078000000078000000078000001FFF80380000000001E000000FC000;
        char[82]     <=  256'h00001E0E070000000038000078078000000FC380300000000001E000007FE000;
        char[83]     <=  256'h00001E060C00000000380003FE07800000000380700000000001C0000FFFC000;
        char[84]     <=  256'h00000E001803C0000038007FFC07800000000380600000000001C007FFFE0000;
        char[85]     <=  256'h00000E0001FFF00000381FFFC007800000000380E00000000001C01FFFC00000;
        char[86]     <=  256'h00000000FFFFFC0000380FF80007800000000380C00000000001CF87E0000000;
        char[87]     <=  256'h0008007FF000FE00003800380003800000000180000F80000001FFC000000000;
        char[88]     <=  256'h000C7FF00001FF000038003C000380000000000007FFE000000FFF8000000000;
        char[89]     <=  256'h001FFC000001FF000038003C0003800000400007FFFFF80001FFFE0000FC0000;
        char[90]     <=  256'h001C00780003C0000038001C0003800000600FFFE003FC000FFFE006007F0000;
        char[91]     <=  256'h003C007C000600000038001C0003800000FFFFC00003FC0003F9C007C03FC000;
        char[92]     <=  256'h0038007C000000000038001CF003800000FFE0F80003F8000003C007C00FC000;
        char[93]     <=  256'h0078007800E000000038001FF803C00001E0007C0007C0000003C007C007E000;
        char[94]     <=  256'h007800781FFC0000003801FFF003C00001E0007C000E00000007C00F8001E000;
        char[95]     <=  256'h00F00073FFF8000000380FFFC003C00003C00078000800000007C01E00000000;
        char[96]     <=  256'h00E000FFFE00000000380FFC0003C00003C0007801C00000000FC03C01C00000;
        char[97]     <=  256'h00E03FFE000000000038003C3803C00007C000383FF00000000FC07001E00000;
        char[98]     <=  256'h0001FFE000000000003800383E03C0000780003FFFF00000001DF8E001F00000;
        char[99]     <=  256'h000001C000000000003800380F03C00007800FFFFFF00000003DFE0001F00000;
        char[100]     <=  256'h000001C000000000003800380703C000070FFFFF800000000039BE1E01E00000;
        char[101]     <=  256'h000003801C000000003000380003C000070FFFF80000000000799E0F01E00000;
        char[102]     <=  256'h00000380FF000000003000380003C0000007C1FC0000000000F18E0783C00000;
        char[103]     <=  256'h000007FFFF800000007000380003C000000003FE0000000001E18003C3C00000;
        char[104]     <=  256'h00000FFE0FC00000007000383F83C000000007B70000000003C38001E7800000;
        char[105]     <=  256'h00000E000F8000000070003FFFE3C00000000F338000000007838000E7800000;
        char[106]     <=  256'h00001FC01F0000000071FFFFFFE3C00000000E31C0000000070380007F000000;
        char[107]     <=  256'h00003CF81E0000000070FF000003C00000001E38E00000000E0380003F000000;
        char[108]     <=  256'h0000783C3C000000007000000003C00000003C38780000001C0380001E000000;
        char[109]     <=  256'h0000701E38000000007000000007C000000078383C000000300380003E000000;
        char[110]     <=  256'h0000E007F8000000007000000007C0000000F0383E000000600380007F000000;
        char[111]     <=  256'h0001C003F000000000F000000007C0000001E0781F80000000038000FFC00000;
        char[112]     <=  256'h00038001F000000000F00001FF87C0000003C0780FE0000000038003F3E00000;
        char[113]     <=  256'h00070003FC00000000F003FFFFC7C000000F807807FC000000078007C1F80000;
        char[114]     <=  256'h000E000FFE00000000FFFFFFFFE7C000001F007803FF80000007801F80FE0000;
        char[115]     <=  256'h001C003E3F80000000FFFE0000FFC000003C007801FFF8000007803E007F8000;
        char[116]     <=  256'h007800FC0FE0000000F00000003FC00000F8007800FFFE00000781F8003FF000;
        char[117]     <=  256'h00E007F007FC000000E00000003F800001E00078007FFC00000F87E0003FFE00;
        char[118]     <=  256'h01C03FC003FFC00000600000001F8000078000F8001F0000000F8000001FFFE0;
        char[119]     <=  256'h0701FC0001FFFE0000600000000F80000C0000F80000000000078000000FFFF0;
        char[120]     <=  256'h00000000007FFFC000000000000F0000000000F800000000000780000007FFE0;
        char[121]     <=  256'h00000000003FFE000000000000070000000000F800000000000700000000F000;
        char[122]     <=  256'h00000000000600000000000000060000000000F8000000000003000000000000;
        char[123]     <=  256'h0000000000000000000000000000000000000078000000000000000000000000;
        char[124]     <=  256'h0000000000000000000000000000000000000070000000000000000000000000;
        char[125]     <=  256'h0000000000000000000000000000000000000000000000000000000000000000;
        char[126]     <=  256'h0000000000000000000000000000000000000000000000000000000000000000;
        char[127]     <=  256'h0000000000000000000000000000000000000000000000000000000000000000;
    end

//pix_data:������ص�ɫ����Ϣ,���ݵ�ǰ���ص�����ָ����ǰ���ص���ɫ����
always@(posedge tft_clk or negedge sys_rst_n)
    if(sys_rst_n == 1'b0)
        pix_data    <= BLACK;
    else    if(((pix_x >= CHAR_B_H) && (pix_x < (CHAR_B_H + CHAR_W)))
                && ((pix_y >= CHAR_B_V) && (pix_y < (CHAR_B_V + CHAR_H))))
        begin
            if(char[char_y][10'd255 - char_x] == 1'b1)
                pix_data    <=  GOLDEN;
            else
                pix_data    <=  BLACK;
        end
    else
        pix_data    <= BLACK;

endmodule